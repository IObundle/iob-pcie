// PCIE

      input PCIE_CLK,
      input PCIE_RST,
      input PCIE_CHNL_RX,
      output PCIE_CHNL_RX_CLK,
      output PCIE_CHNL_RX_ACK,
      input PCIE_CHNL_RX_LAST,
      input [31:0] PCIE_CHNL_RX_LEN,
      input [30:0] PCIE_CHNL_RX_OFF,
      input [31:0] PCIE_CHNL_RX_DATA,
      input PCIE_CHNL_RX_DATA_VALID,
      output PCIE_CHNL_RX_DATA_REN,
      output PCIE_CHNL_TX_CLK,
      output PCIE_CHNL_TX,
      input PCIE_CHNL_TX_ACK,
      output PCIE_CHNL_TX_LAST,
      output [31:0] PCIE_CHNL_TX_LEN,
      output [30:0] PCIE_CHNL_TX_OFF,
      output [31:0] PCIE_CHNL_TX_DATA,
      output PCIE_CHNL_TX_DATA_VALID,
      input PCIE_CHNL_TX_DATA_REN,
